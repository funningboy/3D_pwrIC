module bench_1_L2 (clk1_OUT ,n256_OUT ,n222_OUT ,N1072_OUT ,N6_OUT ,n246_OUT ,n200_OUT ,n255_OUT ,n176_OUT ,n247_OUT ,n216_OUT ,N331_OUT ,n252_OUT ,N4_OUT ,N168_OUT ,N10_OUT ,n249_OUT ,N26_OUT ,N334_OUT ,n234_OUT ,N31_OUT ,N23_OUT ,N6_OUT ,n258_OUT ,n257_OUT ,N4_OUT ,N14_OUT ,n260_OUT ,N106_OUT ,n209_OUT ,n212_OUT ,n253_OUT ,n186_OUT ,n183_OUT ,N331_OUT,n208_IN ,n219_IN ,N27_IN ,n211_IN ,N5_IN ,N168_IN ,n256_IN ,n264_IN ,n231_IN ,N1070_IN ,n199_IN ,N15_IN ,N32_IN ,clk1_IN ,N334_IN ,n243_IN ,N31_IN ,n175_IN ,n171_IN ,N7_IN ,N11_IN ,n249_IN ,N24_IN ,clk2_IN ,n257_IN ,n195_IN ,N25_IN ,n258_IN ,n262_IN ,n254_IN ,X34_IN ,n260_IN ,X0_IN ,n255_IN ,N1071_IN ,N23_IN ,n248_IN);

output clk1_OUT ,n256_OUT ,n222_OUT ,N1072_OUT ,N6_OUT ,n246_OUT ,n200_OUT ,n255_OUT ,n176_OUT ,n247_OUT ,n216_OUT ,N331_OUT ,n252_OUT ,N4_OUT ,N168_OUT ,N10_OUT ,n249_OUT ,N26_OUT ,N334_OUT ,n234_OUT ,N31_OUT ,N23_OUT ,N6_OUT ,n258_OUT ,n257_OUT ,N4_OUT ,N14_OUT ,n260_OUT ,N106_OUT ,n209_OUT ,n212_OUT ,n253_OUT ,n186_OUT ,n183_OUT ,N331_OUT;

input n208_IN ,n219_IN ,N27_IN ,n211_IN ,N5_IN ,N168_IN ,n256_IN ,n264_IN ,n231_IN ,N1070_IN ,n199_IN ,N15_IN ,N32_IN ,clk1_IN ,N334_IN ,n243_IN ,N31_IN ,n175_IN ,n171_IN ,N7_IN ,N11_IN ,n249_IN ,N24_IN ,clk2_IN ,n257_IN ,n195_IN ,N25_IN ,n258_IN ,n262_IN ,n254_IN ,X34_IN ,n260_IN ,X0_IN ,n255_IN ,N1071_IN ,N23_IN ,n248_IN;

AND2X1 U312_ ( .A(N19) , .B(n207) , .Y(n210) );
AND2X1 U308_ ( .B(n219) , .A(N15) , .Y(n222) );
AND2X1 U316_ ( .B(n195) , .A(N23) , .Y(n198) );
AND2X1 U315_ ( .B(n198) , .A(N22) , .Y(n201) );
AND2X1 U304_ ( .A(N11) , .B(n231) , .Y(n234) );
AND2X1 U314_ ( .A(N21) , .B(n201) , .Y(n204) );
AND2X1 U310_ ( .B(n213) , .A(N17) , .Y(n216) );
AND2X1 U313_ ( .B(n204) , .A(N20) , .Y(n207) );
AND2X1 U311_ ( .B(n210) , .A(N18) , .Y(n213) );
AND2X2 U298_ ( .B(n249) , .A(N5) , .Y(n252) );
AND2X2 U103_ ( .B(N1083) , .A(N1071) , .Y(N1082) );
AND2X2 U323_ ( .B(n174) , .A(N30) , .Y(n177) );
AND2X2 U322_ ( .A(N29) , .B(n177) , .Y(n180) );
AND2X2 U321_ ( .B(n180) , .A(N28) , .Y(n183) );
AND2X2 U320_ ( .B(n183) , .A(N27) , .Y(n186) );
AND2X2 U300_ ( .A(N7) , .B(n243) , .Y(n246) );
DFFX1 DFF14_ ( .CK(clk1) , .D(N231) , .Q(N14) );
DFFX1 DFF6_ ( .D(N287) , .CK(clk1) , .Q(N6) );
DFFX1 DFF35_ ( .CK(clk2) , .D(N335) , .Q(N333) );
DFFX1 DFF10_ ( .CK(clk1) , .D(N259) , .Q(N10) );
DFFX1 DFF4_ ( .D(N301) , .CK(clk1) , .Q(N4) );
DFFX1 DFF33_ ( .D(X0) , .CK(clk2) , .Q(N331) );
DFFX2 DFF19_ ( .D(N196) , .CK(clk1) , .Q(N19) );
DFFX2 DFF18_ ( .D(N203) , .CK(clk1) , .Q(N18) );
DFFX2 DFF30_ ( .D(N119) , .CK(clk1) , .Q(N30) );
DFFX2 DFF29_ ( .D(N126) , .CK(clk1) , .Q(N29) );
DFFX2 DFF20_ ( .D(N189) , .CK(clk1) , .Q(N20) );
DFFX2 DFF22_ ( .CK(clk1) , .D(N175) , .Q(N22) );
DFFX2 DFF28_ ( .D(N133) , .CK(clk1) , .Q(N28) );
DFFX2 DFF26_ ( .CK(clk1) , .D(N147) , .Q(N26) );
DFFX2 DFF21_ ( .CK(clk1) , .D(N182) , .Q(N21) );
DFFX2 DFF17_ ( .D(N210) , .CK(clk1) , .Q(N17) );
DFFX2 DFF59_ ( .CK(clk1) , .D(N1082) , .Q(N1072) );
INVX1 U268_ ( .A(N10) , .Y(n233) );
INVX1 U244_ ( .A(N18) , .Y(n209) );
INVX1 U247_ ( .A(N17) , .Y(n212) );
INVX1 U235_ ( .A(N21) , .Y(n200) );
INVX1 U220_ ( .A(N26) , .Y(n185) );
INVX1 U214_ ( .A(N28) , .Y(n179) );
INVX1 U208_ ( .A(N30) , .Y(n173) );
INVX1 U256_ ( .A(N14) , .Y(n221) );
INVX1 U238_ ( .A(N20) , .Y(n203) );
INVX1 U232_ ( .A(N22) , .Y(n197) );
INVX2 U241_ ( .A(N19) , .Y(n206) );
INVX2 U280_ ( .A(N6) , .Y(n245) );
INVX2 U286_ ( .A(N4) , .Y(n251) );
INVX2 U211_ ( .A(N29) , .Y(n176) );
MX2X1 U245_ ( .B(n212) , .S0(n213) , .A(n211) , .Y(N210) );
MX2X1 U209_ ( .S0(n177) , .B(n176) , .A(n175) , .Y(N126) );
MX2X1 U230_ ( .B(n197) , .S0(n198) , .A(n196) , .Y(N175) );
MX2X1 U233_ ( .B(n200) , .S0(n201) , .A(n199) , .Y(N182) );
MX2X1 U254_ ( .S0(n222) , .B(n221) , .A(n220) , .Y(N231) );
MX2X1 U206_ ( .S0(n174) , .B(n173) , .A(n172) , .Y(N119) );
MX2X1 U239_ ( .S0(n207) , .B(n206) , .A(n205) , .Y(N196) );
MX2X1 U236_ ( .B(n203) , .A(n202) , .S0(n204) , .Y(N189) );
MX2X1 U218_ ( .S0(n186) , .A(n184) , .B(n185) , .Y(N147) );
MX2X1 U266_ ( .A(n232) , .B(n233) , .S0(n234) , .Y(N259) );
MX2X2 U212_ ( .A(n178) , .S0(n180) , .B(n179) , .Y(N133) );
MX2X2 U278_ ( .S0(n246) , .B(n245) , .A(n244) , .Y(N287) );
MX2X2 U284_ ( .S0(n252) , .B(n251) , .A(n250) , .Y(N301) );
MX2X2 U242_ ( .B(n209) , .S0(n210) , .A(n208) , .Y(N203) );
NAND4X2 U337_ ( .C(N19) , .B(N18) , .D(N20) , .A(N17) , .Y(n270) );
NAND4X2 U336_ ( .A(N29) , .B(N30) , .D(N32) , .C(N31) , .Y(n271) );
NAND4X2 U335_ ( .B(N26) , .D(N28) , .A(N25) , .C(N27) , .Y(n272) );
NAND4X2 U338_ ( .A(N21) , .B(N22) , .C(N23) , .D(N24) , .Y(n269) );
NOR2X1 U267_ ( .B(n233) , .A(N333) , .Y(n232) );
NOR2X1 U285_ ( .B(n251) , .A(N333) , .Y(n250) );
NOR2X1 U219_ ( .A(N333) , .B(n185) , .Y(n184) );
NOR2X1 U255_ ( .B(n221) , .A(N333) , .Y(n220) );
NOR2X1 U237_ ( .B(n203) , .A(N333) , .Y(n202) );
NOR2X1 U240_ ( .B(n206) , .A(N334) , .Y(n205) );
NOR2X2 U279_ ( .B(n245) , .A(N333) , .Y(n244) );
NOR2X2 U328_ ( .A(n263) , .B(n264) , .Y(N106) );
NOR2X2 U288_ ( .B(n254) , .A(N334) , .Y(n253) );
NOR2X2 U282_ ( .A(N334) , .B(n248) , .Y(n247) );
NOR3X2 U324_ ( .B(N331) , .A(n262) , .C(n171) , .Y(n174) );
OR2X2 U119_ ( .A(X34) , .B(X0) , .Y(N335) );
OR4X2 U334_ ( .D(n272) , .C(n271) , .B(n270) , .A(n269) , .Y(n263) );
TSV_CELL TSV_CELL_63_ ( .DN(n219_IN) , .UP(n219) );
TSV_CELL TSV_CELL_54_ ( .UP(n222) , .DN(n222_OUT) );
TSV_CELL TSV_CELL_21_ ( .UP(N1072) , .DN(N1072_OUT) );
TSV_CELL TSV_CELL_51_ ( .UP(N6) , .DN(N6_OUT) );
TSV_CELL TSV_CELL_26_ ( .DN(N27_IN) , .UP(N27) );
TSV_CELL TSV_CELL_67_ ( .DN(n211_IN) , .UP(n211) );
TSV_CELL TSV_CELL_11_ ( .DN(N5_IN) , .UP(N5) );
TSV_CELL TSV_CELL_57_ ( .UP(n255) , .DN(n255_OUT) );
TSV_CELL TSV_CELL_68_ ( .DN(N168_IN) , .UP(N168) );
TSV_CELL TSV_CELL_59_ ( .UP(n176) , .DN(n176_OUT) );
TSV_CELL TSV_CELL_62_ ( .UP(n247) , .DN(n247_OUT) );
TSV_CELL TSV_CELL_1_ ( .UP(n216) , .DN(n216_OUT) );
TSV_CELL TSV_CELL_40_ ( .DN(n256_IN) , .UP(n256) );
TSV_CELL TSV_CELL_53_ ( .DN(n264_IN) , .UP(n264) );
TSV_CELL TSV_CELL_27_ ( .DN(n231_IN) , .UP(n231) );
TSV_CELL TSV_CELL_4_ ( .DN(N1070_IN) , .UP(N1070) );
TSV_CELL TSV_CELL_55_ ( .DN(N15_IN) , .UP(N15) );
TSV_CELL TSV_CELL_22_ ( .DN(N32_IN) , .UP(N32) );
TSV_CELL TSV_CELL_32_ ( .UP(N10) , .DN(N10_OUT) );
TSV_CELL TSV_CELL_7_ ( .UP(n249) , .DN(n249_OUT) );
TSV_CELL TSV_CELL_30_ ( .DN(clk1_IN) , .UP(clk1) );
TSV_CELL TSV_CELL_46_ ( .DN(N334_IN) , .UP(N334) );
TSV_CELL TSV_CELL_19_ ( .UP(N26) , .DN(N26_OUT) );
TSV_CELL TSV_CELL_60_ ( .DN(n243_IN) , .UP(n243) );
TSV_CELL TSV_CELL_34_ ( .DN(N31_IN) , .UP(N31) );
TSV_CELL TSV_CELL_25_ ( .DN(n175_IN) , .UP(n175) );
TSV_CELL TSV_CELL_17_ ( .DN(n171_IN) , .UP(n171) );
TSV_CELL TSV_CELL_56_ ( .DN(N7_IN) , .UP(N7) );
TSV_CELL TSV_CELL_29_ ( .UP(n234) , .DN(n234_OUT) );
TSV_CELL TSV_CELL_61_ ( .DN(N11_IN) , .UP(N11) );
TSV_CELL TSV_CELL_48_ ( .DN(N24_IN) , .UP(N24) );
TSV_CELL TSV_CELL_15_ ( .DN(clk2_IN) , .UP(clk2) );
TSV_CELL TSV_CELL_9_ ( .DN(n195_IN) , .UP(n195) );
TSV_CELL TSV_CELL_49_ ( .UP(N23) , .DN(N23_OUT) );
TSV_CELL TSV_CELL_45_ ( .DN(N25_IN) , .UP(N25) );
TSV_CELL TSV_CELL_37_ ( .DN(n258_IN) , .UP(n258) );
TSV_CELL TSV_CELL_33_ ( .DN(n254_IN) , .UP(n254) );
TSV_CELL TSV_CELL_23_ ( .DN(X34_IN) , .UP(X34) );
TSV_CELL TSV_CELL_13_ ( .UP(n257) , .DN(n257_OUT) );
TSV_CELL TSV_CELL_70_ ( .UP(N4) , .DN(N4_OUT) );
TSV_CELL TSV_CELL_20_ ( .UP(N14) , .DN(N14_OUT) );
TSV_CELL TSV_CELL_0_ ( .DN(X0_IN) , .UP(X0) );
TSV_CELL TSV_CELL_5_ ( .UP(n260) , .DN(n260_OUT) );
TSV_CELL TSV_CELL_16_ ( .UP(N106) , .DN(N106_OUT) );
TSV_CELL TSV_CELL_24_ ( .UP(n212) , .DN(n212_OUT) );
TSV_CELL TSV_CELL_3_ ( .UP(n253) , .DN(n253_OUT) );
TSV_CELL TSV_CELL_36_ ( .UP(n186) , .DN(n186_OUT) );
TSV_CELL TSV_CELL_12_ ( .UP(n183) , .DN(n183_OUT) );
TSV_CELL TSV_CELL_66_ ( .DN(N1071_IN) , .UP(N1071) );
TSV_CELL TSV_CELL_43_ ( .UP(N331) , .DN(N331_OUT) );
TSV_CELL TSV_CELL_39_ ( .DN(n248_IN) , .UP(n248) );
TSV_LAND TSV_LAND_31_ ( .DN(clk1) , .UP(clk1_OUT) );
TSV_LAND TSV_LAND_28_ ( .UP(n208_IN) , .DN(n208) );
TSV_LAND TSV_LAND_41_ ( .DN(n256) , .UP(n256_OUT) );
TSV_LAND TSV_LAND_2_ ( .DN(n246) , .UP(n246_OUT) );
TSV_LAND TSV_LAND_64_ ( .DN(n200) , .UP(n200_OUT) );
TSV_LAND TSV_LAND_44_ ( .DN(N331) , .UP(N331_OUT) );
TSV_LAND TSV_LAND_18_ ( .DN(n252) , .UP(n252_OUT) );
TSV_LAND TSV_LAND_71_ ( .DN(N4) , .UP(N4_OUT) );
TSV_LAND TSV_LAND_69_ ( .DN(N168) , .UP(N168_OUT) );
TSV_LAND TSV_LAND_65_ ( .UP(n199_IN) , .DN(n199) );
TSV_LAND TSV_LAND_47_ ( .DN(N334) , .UP(N334_OUT) );
TSV_LAND TSV_LAND_35_ ( .DN(N31) , .UP(N31_OUT) );
TSV_LAND TSV_LAND_8_ ( .UP(n249_IN) , .DN(n249) );
TSV_LAND TSV_LAND_14_ ( .UP(n257_IN) , .DN(n257) );
TSV_LAND TSV_LAND_52_ ( .DN(N6) , .UP(N6_OUT) );
TSV_LAND TSV_LAND_42_ ( .UP(n262_IN) , .DN(n262) );
TSV_LAND TSV_LAND_6_ ( .UP(n260_IN) , .DN(n260) );
TSV_LAND TSV_LAND_38_ ( .DN(n258) , .UP(n258_OUT) );
TSV_LAND TSV_LAND_58_ ( .UP(n255_IN) , .DN(n255) );
TSV_LAND TSV_LAND_10_ ( .DN(n209) , .UP(n209_OUT) );
TSV_LAND TSV_LAND_50_ ( .UP(N23_IN) , .DN(N23) );
XNOR2X1 U231_ ( .B(n197) , .A(N333) , .Y(n196) );
XNOR2X1 U207_ ( .A(N333) , .B(n173) , .Y(n172) );
XOR2X2 U213_ ( .B(n179) , .A(N331) , .Y(n178) );
XOR2X2 U102_ ( .B(N1072) , .A(N1070) , .Y(N1083) );
endmodule
