module bench_1_L3 (n255_OUT ,N23_OUT ,n262_OUT ,n199_OUT ,n257_OUT ,n249_OUT ,n208_OUT ,n260_OUT,N6_IN ,n200_IN ,N331_IN ,N4_IN ,N31_IN ,n256_IN ,n246_IN ,N168_IN ,clk1_IN ,n252_IN ,n258_IN ,n209_IN ,N334_IN);

output n255_OUT ,N23_OUT ,n262_OUT ,n199_OUT ,n257_OUT ,n249_OUT ,n208_OUT ,n260_OUT;

input N6_IN ,n200_IN ,N331_IN ,N4_IN ,N31_IN ,n256_IN ,n246_IN ,N168_IN ,clk1_IN ,n252_IN ,n258_IN ,n209_IN ,N334_IN;

AND2X2 U299_ ( .A(N6) , .B(n246) , .Y(n249) );
AND2X2 U297_ ( .A(N4) , .B(n252) , .Y(n255) );
DFFX2 DFF23_ ( .CK(clk1) , .D(N168) , .Q(N23) );
INVX1 U326_ ( .A(N31) , .Y(n262) );
NOR2X2 U243_ ( .B(n209) , .A(N331) , .Y(n208) );
NOR2X2 U291_ ( .A(N331) , .B(n256) , .Y(n257) );
OR2X1 U295_ ( .B(n258) , .A(n256) , .Y(n260) );
TSV_CELL TSV_CELL_52_ ( .DN(N6_IN) , .UP(N6) );
TSV_CELL TSV_CELL_64_ ( .DN(n200_IN) , .UP(n200) );
TSV_CELL TSV_CELL_58_ ( .UP(n255) , .DN(n255_OUT) );
TSV_CELL TSV_CELL_44_ ( .DN(N331_IN) , .UP(N331) );
TSV_CELL TSV_CELL_71_ ( .DN(N4_IN) , .UP(N4) );
TSV_CELL TSV_CELL_35_ ( .DN(N31_IN) , .UP(N31) );
TSV_CELL TSV_CELL_41_ ( .DN(n256_IN) , .UP(n256) );
TSV_CELL TSV_CELL_50_ ( .UP(N23) , .DN(N23_OUT) );
TSV_CELL TSV_CELL_2_ ( .DN(n246_IN) , .UP(n246) );
TSV_CELL TSV_CELL_69_ ( .DN(N168_IN) , .UP(N168) );
TSV_CELL TSV_CELL_31_ ( .DN(clk1_IN) , .UP(clk1) );
TSV_CELL TSV_CELL_18_ ( .DN(n252_IN) , .UP(n252) );
TSV_CELL TSV_CELL_42_ ( .UP(n262) , .DN(n262_OUT) );
TSV_CELL TSV_CELL_38_ ( .DN(n258_IN) , .UP(n258) );
TSV_CELL TSV_CELL_65_ ( .UP(n199) , .DN(n199_OUT) );
TSV_CELL TSV_CELL_10_ ( .DN(n209_IN) , .UP(n209) );
TSV_CELL TSV_CELL_14_ ( .UP(n257) , .DN(n257_OUT) );
TSV_CELL TSV_CELL_8_ ( .UP(n249) , .DN(n249_OUT) );
TSV_CELL TSV_CELL_47_ ( .DN(N334_IN) , .UP(N334) );
TSV_CELL TSV_CELL_28_ ( .UP(n208) , .DN(n208_OUT) );
TSV_CELL TSV_CELL_6_ ( .UP(n260) , .DN(n260_OUT) );
XNOR2X2 U234_ ( .B(n200) , .A(N334) , .Y(n199) );
endmodule
