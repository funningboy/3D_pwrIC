module _ic3d_top_ (X1061,X0 ,X1 ,X34 ,clk1 ,clk2);

output X1061;

input X0 ,X1 ,X34 ,clk1 ,clk2;

bench_1_L0 i_bench_1_L0 ( .X1061_IN(X1061_10) , .clk1_OUT(clk1_01) , .X0_OUT(X0_01) , .X34_OUT(X34_01) , .clk2_OUT(clk2_01) , .X1_OUT(X1_01) );

bench_1_L1 i_bench_1_L1 ( .clk1_IN(clk1_01) , .clk2_IN(clk2_01) , .X1_IN(X1_01) , .N4_IN(N4_21) , .N26_IN(N26_21) , .X34_IN(X34_01) , .n257_IN(n257_21) , .n212_IN(n212_21) , .n255_IN(n255_21) , .N6_IN(N6_21) , .N106_IN(N106_21) , .n253_IN(n253_21) , .N14_IN(N14_21) , .N23_IN(N23_21) , .n216_IN(n216_21) , .n176_IN(n176_21) , .n234_IN(n234_21) , .n249_IN(n249_21) , .n260_IN(n260_21) , .N331_IN(N331_21) , .n247_IN(n247_21) , .n183_IN(n183_21) , .n186_IN(n186_21) , .X0_IN(X0_01) , .N1072_IN(N1072_21) , .n222_IN(n222_21) , .N10_IN(N10_21) , .n195_OUT(n195_12) , .N1071_OUT(N1071_12) , .n254_OUT(n254_12) , .clk2_OUT(clk2_12) , .N27_OUT(N27_12) , .N11_OUT(N11_12) , .X34_OUT(X34_12) , .N15_OUT(N15_12) , .n211_OUT(n211_12) , .n243_OUT(n243_12) , .N168_OUT(N168_12) , .N25_OUT(N25_12) , .N32_OUT(N32_12) , .n231_OUT(n231_12) , .n171_OUT(n171_12) , .n256_OUT(n256_12) , .n264_OUT(n264_12) , .N31_OUT(N31_12) , .N1070_OUT(N1070_12) , .X1061_OUT(X1061_10) , .n175_OUT(n175_12) , .n219_OUT(n219_12) , .N334_OUT(N334_12) , .n248_OUT(n248_12) , .n258_OUT(n258_12) , .N7_OUT(N7_12) , .X0_OUT(X0_12) , .clk1_OUT(clk1_12) , .N5_OUT(N5_12) , .N24_OUT(N24_12) );

bench_1_L2 i_bench_1_L2 ( .n208_IN(n208_32) , .n219_IN(n219_12) , .N27_IN(N27_12) , .n211_IN(n211_12) , .N5_IN(N5_12) , .N168_IN(N168_12) , .n256_IN(n256_12) , .n264_IN(n264_12) , .n231_IN(n231_12) , .N1070_IN(N1070_12) , .n199_IN(n199_32) , .N15_IN(N15_12) , .N32_IN(N32_12) , .clk1_IN(clk1_12) , .N334_IN(N334_12) , .n243_IN(n243_12) , .N31_IN(N31_12) , .n175_IN(n175_12) , .n171_IN(n171_12) , .N7_IN(N7_12) , .N11_IN(N11_12) , .n249_IN(n249_32) , .N24_IN(N24_12) , .clk2_IN(clk2_12) , .n257_IN(n257_32) , .n195_IN(n195_12) , .N25_IN(N25_12) , .n258_IN(n258_12) , .n262_IN(n262_32) , .n254_IN(n254_12) , .X34_IN(X34_12) , .n260_IN(n260_32) , .X0_IN(X0_12) , .n255_IN(n255_32) , .N1071_IN(N1071_12) , .N23_IN(N23_32) , .n248_IN(n248_12) , .clk1_OUT(clk1_23) , .n256_OUT(n256_23) , .n222_OUT(n222_21) , .N1072_OUT(N1072_21) , .N6_OUT(N6_21) , .n246_OUT(n246_23) , .n200_OUT(n200_23) , .n255_OUT(n255_21) , .n176_OUT(n176_21) , .n247_OUT(n247_21) , .n216_OUT(n216_21) , .N331_OUT(N331_23) , .n252_OUT(n252_23) , .N4_OUT(N4_23) , .N168_OUT(N168_23) , .N10_OUT(N10_21) , .n249_OUT(n249_21) , .N26_OUT(N26_21) , .N334_OUT(N334_23) , .n234_OUT(n234_21) , .N31_OUT(N31_23) , .N23_OUT(N23_21) , .N6_OUT(N6_23) , .n258_OUT(n258_23) , .n257_OUT(n257_21) , .N4_OUT(N4_21) , .N14_OUT(N14_21) , .n260_OUT(n260_21) , .N106_OUT(N106_21) , .n209_OUT(n209_23) , .n212_OUT(n212_21) , .n253_OUT(n253_21) , .n186_OUT(n186_21) , .n183_OUT(n183_21) , .N331_OUT(N331_21) );

bench_1_L3 i_bench_1_L3 ( .N6_IN(N6_23) , .n200_IN(n200_23) , .N331_IN(N331_23) , .N4_IN(N4_23) , .N31_IN(N31_23) , .n256_IN(n256_23) , .n246_IN(n246_23) , .N168_IN(N168_23) , .clk1_IN(clk1_23) , .n252_IN(n252_23) , .n258_IN(n258_23) , .n209_IN(n209_23) , .N334_IN(N334_23) , .n255_OUT(n255_32) , .N23_OUT(N23_32) , .n262_OUT(n262_32) , .n199_OUT(n199_32) , .n257_OUT(n257_32) , .n249_OUT(n249_32) , .n208_OUT(n208_32) , .n260_OUT(n260_32) );

endmodule
