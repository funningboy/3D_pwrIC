module bench_1 ( X0, X1, X34, X1061, 
                 clk1, clk2 );
  input X0, X1, X34, clk1, clk2;
  output X1061;
  
  
  DFFX1 DFF1 ( .Q(N1), .D(N320), .CK(clk1) );
  DFFX1 DFF2 ( .Q(N2), .D(N315), .CK(clk1) );
  DFFX1 DFF3 ( .Q(N3), .D(N308), .CK(clk1) );
  DFFX1 DFF4 ( .Q(N4), .D(N301), .CK(clk1) );
  DFFX1 DFF5 ( .Q(N5), .D(N294), .CK(clk1) );
  DFFX1 DFF6 ( .Q(N6), .D(N287), .CK(clk1) );
  DFFX1 DFF7 ( .Q(N7), .D(N280), .CK(clk1) );
  DFFX1 DFF8 ( .Q(N8), .D(N273), .CK(clk1) );
  DFFX1 DFF9 ( .Q(N9), .D(N266), .CK(clk1) );
  DFFX1 DFF10 ( .Q(N10), .D(N259), .CK(clk1) );
  DFFX1 DFF11 ( .Q(N11), .D(N252), .CK(clk1) );
  DFFX1 DFF12 ( .Q(N12), .D(N245), .CK(clk1) );
  DFFX1 DFF13 ( .Q(N13), .D(N238), .CK(clk1) );
  DFFX1 DFF14 ( .Q(N14), .D(N231), .CK(clk1) );
  DFFX1 DFF15 ( .Q(N15), .D(N224), .CK(clk1) );
  DFFX1 DFF16 ( .Q(N16), .D(N217), .CK(clk1) );
  DFFX2 DFF17 ( .Q(N17), .D(N210), .CK(clk1) );
  DFFX2 DFF18 ( .Q(N18), .D(N203), .CK(clk1) );
  DFFX2 DFF19 ( .Q(N19), .D(N196), .CK(clk1) );
  DFFX2 DFF20 ( .Q(N20), .D(N189), .CK(clk1) );
  DFFX2 DFF21 ( .Q(N21), .D(N182), .CK(clk1) );
  DFFX2 DFF22 ( .Q(N22), .D(N175), .CK(clk1) );
  DFFX2 DFF23 ( .Q(N23), .D(N168), .CK(clk1) );
  DFFX2 DFF24 ( .Q(N24), .D(N161), .CK(clk1) );
  DFFX2 DFF25 ( .Q(N25), .D(N154), .CK(clk1) );
  DFFX2 DFF26 ( .Q(N26), .D(N147), .CK(clk1) );
  DFFX2 DFF27 ( .Q(N27), .D(N140), .CK(clk1) );
  DFFX2 DFF28 ( .Q(N28), .D(N133), .CK(clk1) );
  DFFX2 DFF29 ( .Q(N29), .D(N126), .CK(clk1) );
  DFFX2 DFF30 ( .Q(N30), .D(N119), .CK(clk1) );
  DFFX2 DFF31 ( .Q(N31), .D(N112), .CK(clk1) );
  DFFX2 DFF32 ( .Q(N32), .D(N102), .CK(clk1) );

  DFFX1 DFF33 ( .Q(N331), .D(X0), .CK(clk2) );
  DFFX1 DFF34 ( .Q(N332), .D(X1), .CK(clk2) );
  DFFX1 DFF35 ( .Q(N333), .D(N335), .CK(clk2) );
  DFFX1 DFF36 ( .Q(N334), .D(N336), .CK(clk2) );

  DFFX2 DFF41 ( .Q(X1061), .D(N1061), .CK(clk2) );
  DFFX2 DFF42 ( .Q(X1062), .D(N1062), .CK(clk2) );

  DFFX2 DFF57 ( .Q(N1070), .D(N1080), .CK(clk1) );
  DFFX2 DFF58 ( .Q(N1071), .D(N1081), .CK(clk1) );
  DFFX2 DFF59 ( .Q(N1072), .D(N1082), .CK(clk1) );

  NOR2X2 U100 ( .A(N1), .B(N1070), .Y(N1080));
  XOR2X1 U101 ( .A(N1070), .B(N1071), .Y(N1081));
  XOR2X2 U102 ( .A(N1070), .B(N1072), .Y(N1083));
  AND2X2 U103 ( .A(N1071), .B(N1083), .Y(N1082));
  INVX1 U104 ( .A(N1070), .Y(N1090));
  INVX1 U105 ( .A(N1071), .Y(N1091));
  INVX1 U106 ( .A(N1072), .Y(N1092));
  AND4X1 U107 ( .A(N106), .B(N1090), .C(N1091), .D(N1092), .Y(N1051));
  AND4X1 U108 ( .A(N106), .B(N1070), .C(N1091), .D(N1092), .Y(N1052));
  AND4X1 U109 ( .A(N106), .B(N1090), .C(N1071), .D(N1092), .Y(N1053));
  AND4X1 U110 ( .A(N106), .B(N1070), .C(N1071), .D(N1092), .Y(N1054));
  AND4X1 U111 ( .A(N106), .B(N1090), .C(N1091), .D(N1072), .Y(N1055));
  AND4X1 U112 ( .A(N106), .B(N1070), .C(N1091), .D(N1072), .Y(N1056));
  AND4X1 U113 ( .A(N106), .B(N1090), .C(N1071), .D(N1072), .Y(N1057));
  AND4X1 U114 ( .A(N106), .B(N1070), .C(N1071), .D(N1072), .Y(N1058));
  AND2X1 U115 ( .A(N1051), .B(N1052), .Y(N1065));
  AND2X1 U116 ( .A(N1053), .B(N1054), .Y(N1066));
  AND2X1 U117 ( .A(N1055), .B(N1056), .Y(N1063));
  AND2X1 U118 ( .A(N1057), .B(N1058), .Y(N1064));
  OR2X2 U119 ( .A(X34), .B(X0), .Y(N335));
  OR2X2 U120 ( .A(X34), .B(X1), .Y(N336));
  NOR2X1 U121 ( .A(N1065), .B(N1063), .Y(N1061));
  NOR2X2 U122 ( .A(N1066), .B(N1064), .Y(N1062));

  NOR2X1 U202 ( .A(N331), .B(n169), .Y(N102) );
  XNOR2X2 U203 ( .A(N32), .B(X34), .Y(n169) );
  NOR2X1 U204 ( .A(N332), .B(n170), .Y(N112) );
  XOR2X1 U205 ( .A(n171), .B(N31), .Y(n170) );
  MX2X1 U206 ( .S0(n174), .B(n173), .A(n172), .Y(N119) );
  XNOR2X1 U207 ( .A(N333), .B(n173), .Y(n172) );
  INVX1 U208 ( .A(N30), .Y(n173) );
  MX2X1 U209 ( .S0(n177), .B(n176), .A(n175), .Y(N126) );
  XNOR2X2 U210 ( .A(N334), .B(n176), .Y(n175) );
  INVX2 U211 ( .A(N29), .Y(n176) );
  MX2X2 U212 ( .S0(n180), .B(n179), .A(n178), .Y(N133) );
  XOR2X2 U213 ( .A(N331), .B(n179), .Y(n178) );
  INVX1 U214 ( .A(N28), .Y(n179) );
  MX2X1 U215 ( .S0(n183), .B(n182), .A(n181), .Y(N140) );
  NOR2X1 U216 ( .A(N332), .B(n182), .Y(n181) );
  INVX1 U217 ( .A(N27), .Y(n182) );
  MX2X1 U218 ( .S0(n186), .B(n185), .A(n184), .Y(N147) );
  NOR2X1 U219 ( .A(N333), .B(n185), .Y(n184) );
  INVX1 U220 ( .A(N26), .Y(n185) );
  MX2X1 U221 ( .S0(n189), .B(n188), .A(n187), .Y(N154) );
  XOR2X1 U222 ( .A(N334), .B(n188), .Y(n187) );
  INVX1 U223 ( .A(N25), .Y(n188) );
  MX2X1 U224 ( .S0(n192), .B(n191), .A(n190), .Y(N161) );
  XOR2X1 U225 ( .A(N331), .B(n191), .Y(n190) );
  INVX1 U226 ( .A(N24), .Y(n191) );
  MX2X1 U227 ( .S0(n195), .B(n194), .A(n193), .Y(N168) );
  XNOR2X1 U228 ( .A(N332), .B(n194), .Y(n193) );
  INVX1 U229 ( .A(N23), .Y(n194) );
  MX2X1 U230 ( .S0(n198), .B(n197), .A(n196), .Y(N175) );
  XNOR2X1 U231 ( .A(N333), .B(n197), .Y(n196) );
  INVX1 U232 ( .A(N22), .Y(n197) );
  MX2X1 U233 ( .S0(n201), .B(n200), .A(n199), .Y(N182) );
  XNOR2X2 U234 ( .A(N334), .B(n200), .Y(n199) );
  INVX1 U235 ( .A(N21), .Y(n200) );
  MX2X1 U236 ( .S0(n204), .B(n203), .A(n202), .Y(N189) );
  NOR2X1 U237 ( .A(N333), .B(n203), .Y(n202) );
  INVX1 U238 ( .A(N20), .Y(n203) );
  MX2X1 U239 ( .S0(n207), .B(n206), .A(n205), .Y(N196) );
  NOR2X1 U240 ( .A(N334), .B(n206), .Y(n205) );
  INVX2 U241 ( .A(N19), .Y(n206) );
  MX2X2 U242 ( .S0(n210), .B(n209), .A(n208), .Y(N203) );
  NOR2X2 U243 ( .A(N331), .B(n209), .Y(n208) );
  INVX1 U244 ( .A(N18), .Y(n209) );
  MX2X1 U245 ( .S0(n213), .B(n212), .A(n211), .Y(N210) );
  NOR2X1 U246 ( .A(N332), .B(n212), .Y(n211) );
  INVX1 U247 ( .A(N17), .Y(n212) );
  MX2X1 U248 ( .S0(n216), .B(n215), .A(n214), .Y(N217) );
  XOR2X1 U249 ( .A(N331), .B(n215), .Y(n214) );
  INVX1 U250 ( .A(N16), .Y(n215) );
  MX2X1 U251 ( .S0(n219), .B(n218), .A(n217), .Y(N224) );
  XOR2X1 U252 ( .A(N332), .B(n218), .Y(n217) );
  INVX1 U253 ( .A(N15), .Y(n218) );
  MX2X1 U254 ( .S0(n222), .B(n221), .A(n220), .Y(N231) );
  NOR2X1 U255 ( .A(N333), .B(n221), .Y(n220) );
  INVX1 U256 ( .A(N14), .Y(n221) );
  MX2X1 U257 ( .S0(n225), .B(n224), .A(n223), .Y(N238) );
  NOR2X1 U258 ( .A(N334), .B(n224), .Y(n223) );
  INVX1 U259 ( .A(N13), .Y(n224) );
  MX2X1 U260 ( .S0(n228), .B(n227), .A(n226), .Y(N245) );
  NOR2X1 U261 ( .A(N331), .B(n227), .Y(n226) );
  INVX1 U262 ( .A(N12), .Y(n227) );
  MX2X1 U263 ( .S0(n231), .B(n230), .A(n229), .Y(N252) );
  NOR2X1 U264 ( .A(N332), .B(n230), .Y(n229) );
  INVX1 U265 ( .A(N11), .Y(n230) );
  MX2X1 U266 ( .S0(n234), .B(n233), .A(n232), .Y(N259) );
  NOR2X1 U267 ( .A(N333), .B(n233), .Y(n232) );
  INVX1 U268 ( .A(N10), .Y(n233) );
  MX2X1 U269 ( .S0(n237), .B(n236), .A(n235), .Y(N266) );
  NOR2X1 U270 ( .A(N334), .B(n236), .Y(n235) );
  INVX1 U271 ( .A(N9), .Y(n236) );
  MX2X1 U272 ( .S0(n240), .B(n239), .A(n238), .Y(N273) );
  NOR2X1 U273 ( .A(N331), .B(n239), .Y(n238) );
  INVX1 U274 ( .A(N8), .Y(n239) );
  MX2X1 U275 ( .S0(n243), .B(n242), .A(n241), .Y(N280) );
  NOR2X1 U276 ( .A(N332), .B(n242), .Y(n241) );
  INVX1 U277 ( .A(N7), .Y(n242) );
  MX2X2 U278 ( .S0(n246), .B(n245), .A(n244), .Y(N287) );
  NOR2X2 U279 ( .A(N333), .B(n245), .Y(n244) );
  INVX2 U280 ( .A(N6), .Y(n245) );
  MX2X2 U281 ( .S0(n249), .B(n248), .A(n247), .Y(N294) );
  NOR2X2 U282 ( .A(N334), .B(n248), .Y(n247) );
  INVX2 U283 ( .A(N5), .Y(n248) );
  MX2X2 U284 ( .S0(n252), .B(n251), .A(n250), .Y(N301) );
  NOR2X1 U285 ( .A(N333), .B(n251), .Y(n250) );
  INVX2 U286 ( .A(N4), .Y(n251) );
  MX2X2 U287 ( .S0(n255), .B(n254), .A(n253), .Y(N308) );
  NOR2X2 U288 ( .A(N334), .B(n254), .Y(n253) );
  INVX2 U289 ( .A(N3), .Y(n254) );
  MX2X1 U290 ( .S0(n258), .B(n257), .A(n256), .Y(N315) );
  NOR2X2 U291 ( .A(N331), .B(n256), .Y(n257) );
  NOR2X2 U292 ( .A(N332), .B(n259), .Y(N320) );
  MX2X2 U293 ( .S0(N1), .B(n261), .A(n260), .Y(n259) );
  NOR2X2 U294 ( .A(n258), .B(n256), .Y(n261) );
  OR2X1 U295 ( .A(n256), .B(n258), .Y(n260) );
  NAND2X1 U296 ( .A(N3), .B(n255), .Y(n258) );
  AND2X2 U297 ( .A(N4), .B(n252), .Y(n255) );
  AND2X2 U298 ( .A(N5), .B(n249), .Y(n252) );
  AND2X2 U299 ( .A(N6), .B(n246), .Y(n249) );
  AND2X2 U300 ( .A(N7), .B(n243), .Y(n246) );
  AND2X1 U301 ( .A(N8), .B(n240), .Y(n243) );
  AND2X1 U302 ( .A(N9), .B(n237), .Y(n240) );
  AND2X1 U303 ( .A(N10), .B(n234), .Y(n237) );
  AND2X1 U304 ( .A(N11), .B(n231), .Y(n234) );
  AND2X1 U305 ( .A(N12), .B(n228), .Y(n231) );
  AND2X1 U306 ( .A(N13), .B(n225), .Y(n228) );
  AND2X1 U307 ( .A(N14), .B(n222), .Y(n225) );
  AND2X1 U308 ( .A(N15), .B(n219), .Y(n222) );
  AND2X1 U309 ( .A(N16), .B(n216), .Y(n219) );
  AND2X1 U310 ( .A(N17), .B(n213), .Y(n216) );
  AND2X1 U311 ( .A(N18), .B(n210), .Y(n213) );
  AND2X1 U312 ( .A(N19), .B(n207), .Y(n210) );
  AND2X1 U313 ( .A(N20), .B(n204), .Y(n207) );
  AND2X1 U314 ( .A(N21), .B(n201), .Y(n204) );
  AND2X1 U315 ( .A(N22), .B(n198), .Y(n201) );
  AND2X1 U316 ( .A(N23), .B(n195), .Y(n198) );
  AND2X2 U317 ( .A(N24), .B(n192), .Y(n195) );
  AND2X2 U318 ( .A(N25), .B(n189), .Y(n192) );
  AND2X2 U319 ( .A(N26), .B(n186), .Y(n189) );
  AND2X2 U320 ( .A(N27), .B(n183), .Y(n186) );
  AND2X2 U321 ( .A(N28), .B(n180), .Y(n183) );
  AND2X2 U322 ( .A(N29), .B(n177), .Y(n180) );
  AND2X2 U323 ( .A(N30), .B(n174), .Y(n177) );
  NOR3X2 U324 ( .A(n262), .B(N331), .C(n171), .Y(n174) );
  NAND2X2 U325 ( .A(N32), .B(X34), .Y(n171) );
  INVX1 U326 ( .A(N31), .Y(n262) );
  INVX2 U327 ( .A(N2), .Y(n256) );
  NOR2X2 U328 ( .A(n263), .B(n264), .Y(N106) );
  OR4X1 U329 ( .A(n265), .B(n266), .C(n267), .D(n268), .Y(n264) );
  NAND4X1 U330 ( .A(N9), .B(N10), .C(N11), .D(N12), .Y(n268) );
  NAND4X1 U331 ( .A(N13), .B(N14), .C(N15), .D(N16), .Y(n267) );
  NAND4X1 U332 ( .A(N1), .B(N2), .C(N3), .D(N4), .Y(n266) );
  NAND4X1 U333 ( .A(N5), .B(N6), .C(N7), .D(N8), .Y(n265) );
  OR4X2 U334 ( .A(n269), .B(n270), .C(n271), .D(n272), .Y(n263) );
  NAND4X2 U335 ( .A(N25), .B(N26), .C(N27), .D(N28), .Y(n272) );
  NAND4X2 U336 ( .A(N29), .B(N30), .C(N31), .D(N32), .Y(n271) );
  NAND4X2 U337 ( .A(N17), .B(N18), .C(N19), .D(N20), .Y(n270) );
  NAND4X2 U338 ( .A(N21), .B(N22), .C(N23), .D(N24), .Y(n269) );
endmodule

