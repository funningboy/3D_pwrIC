module bench_1_L1 (n195_OUT ,N1071_OUT ,n254_OUT ,clk2_OUT ,N27_OUT ,N11_OUT ,X34_OUT ,N15_OUT ,n211_OUT ,n243_OUT ,N168_OUT ,N25_OUT ,N32_OUT ,n231_OUT ,n171_OUT ,n256_OUT ,n264_OUT ,N31_OUT ,N1070_OUT ,X1061_OUT ,n175_OUT ,n219_OUT ,N334_OUT ,n248_OUT ,n258_OUT ,N7_OUT ,X0_OUT ,clk1_OUT ,N5_OUT ,N24_OUT,clk1_IN ,clk2_IN ,X1_IN ,N4_IN ,N26_IN ,X34_IN ,n257_IN ,n212_IN ,n255_IN ,N6_IN ,N106_IN ,n253_IN ,N14_IN ,N23_IN ,n216_IN ,n176_IN ,n234_IN ,n249_IN ,n260_IN ,N331_IN ,n247_IN ,n183_IN ,n186_IN ,X0_IN ,N1072_IN ,n222_IN ,N10_IN);

output n195_OUT ,N1071_OUT ,n254_OUT ,clk2_OUT ,N27_OUT ,N11_OUT ,X34_OUT ,N15_OUT ,n211_OUT ,n243_OUT ,N168_OUT ,N25_OUT ,N32_OUT ,n231_OUT ,n171_OUT ,n256_OUT ,n264_OUT ,N31_OUT ,N1070_OUT ,X1061_OUT ,n175_OUT ,n219_OUT ,N334_OUT ,n248_OUT ,n258_OUT ,N7_OUT ,X0_OUT ,clk1_OUT ,N5_OUT ,N24_OUT;

input clk1_IN ,clk2_IN ,X1_IN ,N4_IN ,N26_IN ,X34_IN ,n257_IN ,n212_IN ,n255_IN ,N6_IN ,N106_IN ,n253_IN ,N14_IN ,N23_IN ,n216_IN ,n176_IN ,n234_IN ,n249_IN ,n260_IN ,N331_IN ,n247_IN ,n183_IN ,n186_IN ,X0_IN ,N1072_IN ,n222_IN ,N10_IN;

AND2X1 U118_ ( .B(N1058) , .A(N1057) , .Y(N1064) );
AND2X1 U305_ ( .A(N12) , .B(n228) , .Y(n231) );
AND2X1 U303_ ( .A(N10) , .B(n234) , .Y(n237) );
AND2X1 U301_ ( .B(n240) , .A(N8) , .Y(n243) );
AND2X1 U116_ ( .B(N1054) , .A(N1053) , .Y(N1066) );
AND2X1 U302_ ( .A(N9) , .B(n237) , .Y(n240) );
AND2X1 U117_ ( .A(N1055) , .B(N1056) , .Y(N1063) );
AND2X1 U306_ ( .B(n225) , .A(N13) , .Y(n228) );
AND2X1 U309_ ( .A(N16) , .B(n216) , .Y(n219) );
AND2X1 U115_ ( .B(N1052) , .A(N1051) , .Y(N1065) );
AND2X1 U307_ ( .A(N14) , .B(n222) , .Y(n225) );
AND2X2 U318_ ( .B(n189) , .A(N25) , .Y(n192) );
AND2X2 U317_ ( .B(n192) , .A(N24) , .Y(n195) );
AND2X2 U319_ ( .A(N26) , .B(n186) , .Y(n189) );
AND4X1 U112_ ( .B(N1070) , .D(N1072) , .A(N106) , .C(N1091) , .Y(N1056) );
AND4X1 U109_ ( .A(N106) , .D(N1092) , .B(N1090) , .C(N1071) , .Y(N1053) );
AND4X1 U111_ ( .D(N1072) , .C(N1091) , .B(N1090) , .A(N106) , .Y(N1055) );
AND4X1 U114_ ( .A(N106) , .D(N1072) , .B(N1070) , .C(N1071) , .Y(N1058) );
AND4X1 U110_ ( .A(N106) , .C(N1071) , .B(N1070) , .D(N1092) , .Y(N1054) );
AND4X1 U107_ ( .B(N1090) , .A(N106) , .D(N1092) , .C(N1091) , .Y(N1051) );
AND4X1 U108_ ( .D(N1092) , .C(N1091) , .B(N1070) , .A(N106) , .Y(N1052) );
AND4X1 U113_ ( .C(N1071) , .D(N1072) , .A(N106) , .B(N1090) , .Y(N1057) );
DFFX1 DFF3_ ( .CK(clk1_IN) , .D(N308) , .Q(N3) );
DFFX1 DFF5_ ( .D(N294) , .CK(clk1_IN) , .Q(N5) );
DFFX1 DFF34_ ( .D(X1_IN) , .CK(clk2_IN) , .Q(N332) );
DFFX1 DFF11_ ( .D(N252) , .CK(clk1_IN) , .Q(N11) );
DFFX1 DFF2_ ( .D(N315) , .CK(clk1_IN) , .Q(N2) );
DFFX1 DFF16_ ( .CK(clk1_IN) , .D(N217) , .Q(N16) );
DFFX1 DFF9_ ( .CK(clk1_IN) , .D(N266) , .Q(N9) );
DFFX1 DFF15_ ( .D(N224) , .CK(clk1_IN) , .Q(N15) );
DFFX1 DFF12_ ( .CK(clk1_IN) , .D(N245) , .Q(N12) );
DFFX1 DFF8_ ( .CK(clk1_IN) , .D(N273) , .Q(N8) );
DFFX1 DFF1_ ( .D(N320) , .CK(clk1_IN) , .Q(N1) );
DFFX1 DFF13_ ( .D(N238) , .CK(clk1_IN) , .Q(N13) );
DFFX1 DFF7_ ( .D(N280) , .CK(clk1_IN) , .Q(N7) );
DFFX1 DFF36_ ( .D(N336) , .CK(clk2_IN) , .Q(N334) );
DFFX2 DFF24_ ( .D(N161) , .CK(clk1_IN) , .Q(N24) );
DFFX2 DFF27_ ( .D(N140) , .CK(clk1_IN) , .Q(N27) );
DFFX2 DFF32_ ( .D(N102) , .CK(clk1_IN) , .Q(N32) );
DFFX2 DFF25_ ( .CK(clk1_IN) , .D(N154) , .Q(N25) );
DFFX2 DFF42_ ( .D(N1062) , .CK(clk2_IN) );
DFFX2 DFF57_ ( .CK(clk1_IN) , .D(N1080) , .Q(N1070) );
DFFX2 DFF31_ ( .D(N112) , .CK(clk1_IN) , .Q(N31) );
DFFX2 DFF41_ ( .CK(clk2_IN) , .D(N1061) , .Q(X1061_OUT) );
DFFX2 DFF58_ ( .D(N1081) , .CK(clk1_IN) , .Q(N1071) );
INVX1 U105_ ( .A(N1071) , .Y(N1091) );
INVX1 U253_ ( .A(N15) , .Y(n218) );
INVX1 U250_ ( .A(N16) , .Y(n215) );
INVX1 U223_ ( .A(N25) , .Y(n188) );
INVX1 U271_ ( .A(N9) , .Y(n236) );
INVX1 U274_ ( .A(N8) , .Y(n239) );
INVX1 U277_ ( .A(N7) , .Y(n242) );
INVX1 U104_ ( .A(N1070) , .Y(N1090) );
INVX1 U262_ ( .A(N12) , .Y(n227) );
INVX1 U217_ ( .A(N27) , .Y(n182) );
INVX1 U226_ ( .A(N24) , .Y(n191) );
INVX1 U106_ ( .A(N1072) , .Y(N1092) );
INVX1 U229_ ( .A(N23) , .Y(n194) );
INVX1 U259_ ( .A(N13) , .Y(n224) );
INVX1 U265_ ( .A(N11) , .Y(n230) );
INVX2 U283_ ( .A(N5) , .Y(n248) );
INVX2 U327_ ( .A(N2) , .Y(n256) );
INVX2 U289_ ( .A(N3) , .Y(n254) );
MX2X1 U257_ ( .B(n224) , .S0(n225) , .A(n223) , .Y(N238) );
MX2X1 U263_ ( .B(n230) , .S0(n231) , .A(n229) , .Y(N252) );
MX2X1 U227_ ( .A(n193) , .B(n194) , .S0(n195) , .Y(N168) );
MX2X1 U224_ ( .B(n191) , .S0(n192) , .A(n190) , .Y(N161) );
MX2X1 U248_ ( .S0(n216) , .B(n215) , .A(n214) , .Y(N217) );
MX2X1 U290_ ( .A(n256) , .S0(n258) , .B(n257) , .Y(N315) );
MX2X1 U221_ ( .B(n188) , .A(n187) , .S0(n189) , .Y(N154) );
MX2X1 U260_ ( .A(n226) , .S0(n228) , .B(n227) , .Y(N245) );
MX2X1 U275_ ( .S0(n243) , .A(n241) , .B(n242) , .Y(N280) );
MX2X1 U269_ ( .B(n236) , .A(n235) , .S0(n237) , .Y(N266) );
MX2X1 U215_ ( .A(n181) , .B(n182) , .S0(n183) , .Y(N140) );
MX2X1 U251_ ( .A(n217) , .B(n218) , .S0(n219) , .Y(N224) );
MX2X1 U272_ ( .S0(n240) , .B(n239) , .A(n238) , .Y(N273) );
MX2X2 U281_ ( .S0(n249) , .B(n248) , .A(n247) , .Y(N294) );
MX2X2 U287_ ( .B(n254) , .S0(n255) , .A(n253) , .Y(N308) );
MX2X2 U293_ ( .A(n260) , .B(n261) , .S0(N1) , .Y(n259) );
NAND2X1 U296_ ( .A(N3) , .B(n255) , .Y(n258) );
NAND2X2 U325_ ( .A(N32) , .B(X34_IN) , .Y(n171) );
NAND4X1 U331_ ( .D(N16) , .A(N13) , .B(N14) , .C(N15) , .Y(n267) );
NAND4X1 U333_ ( .C(N7) , .D(N8) , .A(N5) , .B(N6) , .Y(n265) );
NAND4X1 U330_ ( .B(N10) , .A(N9) , .D(N12) , .C(N11) , .Y(n268) );
NAND4X1 U332_ ( .D(N4) , .A(N1) , .B(N2) , .C(N3) , .Y(n266) );
NOR2X1 U273_ ( .B(n239) , .A(N331) , .Y(n238) );
NOR2X1 U261_ ( .A(N331) , .B(n227) , .Y(n226) );
NOR2X1 U264_ ( .A(N332) , .B(n230) , .Y(n229) );
NOR2X1 U204_ ( .A(N332) , .B(n170) , .Y(N112) );
NOR2X1 U276_ ( .B(n242) , .A(N332) , .Y(n241) );
NOR2X1 U270_ ( .A(N334) , .B(n236) , .Y(n235) );
NOR2X1 U246_ ( .B(n212) , .A(N332) , .Y(n211) );
NOR2X1 U202_ ( .A(N331) , .B(n169) , .Y(N102) );
NOR2X1 U258_ ( .B(n224) , .A(N334) , .Y(n223) );
NOR2X1 U121_ ( .A(N1065) , .B(N1063) , .Y(N1061) );
NOR2X1 U216_ ( .A(N332) , .B(n182) , .Y(n181) );
NOR2X2 U100_ ( .B(N1070) , .A(N1) , .Y(N1080) );
NOR2X2 U292_ ( .A(N332) , .B(n259) , .Y(N320) );
NOR2X2 U122_ ( .B(N1064) , .A(N1066) , .Y(N1062) );
NOR2X2 U294_ ( .B(n256) , .A(n258) , .Y(n261) );
OR2X2 U120_ ( .B(X1_IN) , .A(X34_IN) , .Y(N336) );
OR4X1 U329_ ( .C(n267) , .D(n268) , .A(n265) , .B(n266) , .Y(n264) );
TSV_LAND TSV_LAND_9_ ( .DN(n195) , .UP(n195_OUT) );
TSV_LAND TSV_LAND_66_ ( .DN(N1071) , .UP(N1071_OUT) );
TSV_LAND TSV_LAND_33_ ( .DN(n254) , .UP(n254_OUT) );
TSV_LAND TSV_LAND_15_ ( .DN(clk2_IN) , .UP(clk2_OUT) );
TSV_LAND TSV_LAND_26_ ( .DN(N27) , .UP(N27_OUT) );
TSV_LAND TSV_LAND_70_ ( .UP(N4_IN) , .DN(N4) );
TSV_LAND TSV_LAND_19_ ( .UP(N26_IN) , .DN(N26) );
TSV_LAND TSV_LAND_61_ ( .DN(N11) , .UP(N11_OUT) );
TSV_LAND TSV_LAND_23_ ( .DN(X34_IN) , .UP(X34_OUT) );
TSV_LAND TSV_LAND_13_ ( .UP(n257_IN) , .DN(n257) );
TSV_LAND TSV_LAND_55_ ( .DN(N15) , .UP(N15_OUT) );
TSV_LAND TSV_LAND_67_ ( .DN(n211) , .UP(n211_OUT) );
TSV_LAND TSV_LAND_60_ ( .DN(n243) , .UP(n243_OUT) );
TSV_LAND TSV_LAND_24_ ( .UP(n212_IN) , .DN(n212) );
TSV_LAND TSV_LAND_68_ ( .DN(N168) , .UP(N168_OUT) );
TSV_LAND TSV_LAND_45_ ( .DN(N25) , .UP(N25_OUT) );
TSV_LAND TSV_LAND_22_ ( .DN(N32) , .UP(N32_OUT) );
TSV_LAND TSV_LAND_57_ ( .UP(n255_IN) , .DN(n255) );
TSV_LAND TSV_LAND_51_ ( .UP(N6_IN) , .DN(N6) );
TSV_LAND TSV_LAND_16_ ( .UP(N106_IN) , .DN(N106) );
TSV_LAND TSV_LAND_27_ ( .DN(n231) , .UP(n231_OUT) );
TSV_LAND TSV_LAND_3_ ( .UP(n253_IN) , .DN(n253) );
TSV_LAND TSV_LAND_17_ ( .DN(n171) , .UP(n171_OUT) );
TSV_LAND TSV_LAND_40_ ( .DN(n256) , .UP(n256_OUT) );
TSV_LAND TSV_LAND_53_ ( .DN(n264) , .UP(n264_OUT) );
TSV_LAND TSV_LAND_20_ ( .UP(N14_IN) , .DN(N14) );
TSV_LAND TSV_LAND_34_ ( .DN(N31) , .UP(N31_OUT) );
TSV_LAND TSV_LAND_49_ ( .UP(N23_IN) , .DN(N23) );
TSV_LAND TSV_LAND_4_ ( .DN(N1070) , .UP(N1070_OUT) );
TSV_LAND TSV_LAND_1_ ( .UP(n216_IN) , .DN(n216) );
TSV_LAND TSV_LAND_59_ ( .UP(n176_IN) , .DN(n176) );
TSV_LAND TSV_LAND_25_ ( .DN(n175) , .UP(n175_OUT) );
TSV_LAND TSV_LAND_29_ ( .UP(n234_IN) , .DN(n234) );
TSV_LAND TSV_LAND_63_ ( .DN(n219) , .UP(n219_OUT) );
TSV_LAND TSV_LAND_46_ ( .DN(N334) , .UP(N334_OUT) );
TSV_LAND TSV_LAND_7_ ( .UP(n249_IN) , .DN(n249) );
TSV_LAND TSV_LAND_39_ ( .DN(n248) , .UP(n248_OUT) );
TSV_LAND TSV_LAND_5_ ( .UP(n260_IN) , .DN(n260) );
TSV_LAND TSV_LAND_43_ ( .UP(N331_IN) , .DN(N331) );
TSV_LAND TSV_LAND_37_ ( .DN(n258) , .UP(n258_OUT) );
TSV_LAND TSV_LAND_62_ ( .UP(n247_IN) , .DN(n247) );
TSV_LAND TSV_LAND_12_ ( .UP(n183_IN) , .DN(n183) );
TSV_LAND TSV_LAND_56_ ( .DN(N7) , .UP(N7_OUT) );
TSV_LAND TSV_LAND_36_ ( .UP(n186_IN) , .DN(n186) );
TSV_LAND TSV_LAND_0_ ( .DN(X0_IN) , .UP(X0_OUT) );
TSV_LAND TSV_LAND_30_ ( .DN(clk1_IN) , .UP(clk1_OUT) );
TSV_LAND TSV_LAND_21_ ( .UP(N1072_IN) , .DN(N1072) );
TSV_LAND TSV_LAND_54_ ( .UP(n222_IN) , .DN(n222) );
TSV_LAND TSV_LAND_11_ ( .DN(N5) , .UP(N5_OUT) );
TSV_LAND TSV_LAND_48_ ( .DN(N24) , .UP(N24_OUT) );
TSV_LAND TSV_LAND_32_ ( .UP(N10_IN) , .DN(N10) );
XNOR2X1 U228_ ( .B(n194) , .A(N332) , .Y(n193) );
XNOR2X2 U210_ ( .B(n176) , .A(N334) , .Y(n175) );
XNOR2X2 U203_ ( .A(N32) , .B(X34_IN) , .Y(n169) );
XOR2X1 U205_ ( .A(n171) , .B(N31) , .Y(n170) );
XOR2X1 U252_ ( .A(N332) , .B(n218) , .Y(n217) );
XOR2X1 U225_ ( .A(N331) , .B(n191) , .Y(n190) );
XOR2X1 U101_ ( .B(N1071) , .A(N1070) , .Y(N1081) );
XOR2X1 U249_ ( .B(n215) , .A(N331) , .Y(n214) );
XOR2X1 U222_ ( .B(n188) , .A(N334) , .Y(n187) );
endmodule
